//interface
interface fs_if;
logic a;
logic b;
logic bin;
logic difference;
logic borrow;
endinterface

//interface.sv
interface fulladder_if;
  logic A;
  logic B;
  logic Cin;
  logic SUM;
  logic CARRY;
endinterface

//transaction.sv
class transaction;
  randc bit A;
  randc bit B;
  randc bit Cin;
  bit SUM ;
  bit CARRY;
endclass

//transaction.sv
class transaction;
  
randc bit a;
randc bit b; 

bit borrow;
bit difference;
  
endclass

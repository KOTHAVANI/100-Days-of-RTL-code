//transaction.sv
class transaction;
randc bit a;
randc bit b;
randc bit bin; 
bit difference;
bit borrow;
endclass

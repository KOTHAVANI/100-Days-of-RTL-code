//interface
interface Seven_Segment_Display_if;
  
  logic [3:0] bcd;
  logic [7:0] segment;

endinterface

//interface
interface transmissiongate_if;
  
  logic  a;
  logic  control;  
  logic  y;
 
endinterface

//interface
interface par_gen_if;
  
logic x;
logic y;
logic z;
logic result;
  
endinterface

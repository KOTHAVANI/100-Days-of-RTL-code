//transaction.sv
class transaction;
  
randc bit x;
randc bit y; 
randc bit z;
bit result;
  
endclass

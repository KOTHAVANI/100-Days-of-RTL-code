//transaction.sv
class transaction;
  
  randc bit [3:0] bcd;
  bit[7:0] segment ;

endclass

//interface
interface hs_if;
  
logic a;
logic b;
logic borrow;
logic difference;
  
endinterface

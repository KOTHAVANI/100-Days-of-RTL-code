`timescale 1ps/1ps
module clock_freq(clock);
input clock;
endmodule

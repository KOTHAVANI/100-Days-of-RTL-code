//transaction.sv
class transaction;
  randc bit a ;
  randc bit control;
   bit  y;
endclass
